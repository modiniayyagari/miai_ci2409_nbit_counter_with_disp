VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter_top
  CLASS BLOCK ;
  FOREIGN counter_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END clk
  PIN cnt_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2099.530 1756.000 2099.810 1760.000 ;
    END
  END cnt_rst
  PIN cnt_start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 233.770 1756.000 234.050 1760.000 ;
    END
  END cnt_start
  PIN cnt_stop
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1166.650 1756.000 1166.930 1760.000 ;
    END
  END cnt_stop
  PIN disp_val[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END disp_val[0]
  PIN disp_val[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1347.800 4.000 1348.400 ;
    END
  END disp_val[10]
  PIN disp_val[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.920 4.000 1473.520 ;
    END
  END disp_val[11]
  PIN disp_val[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1598.040 4.000 1598.640 ;
    END
  END disp_val[12]
  PIN disp_val[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.160 4.000 1723.760 ;
    END
  END disp_val[13]
  PIN disp_val[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END disp_val[1]
  PIN disp_val[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END disp_val[2]
  PIN disp_val[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END disp_val[3]
  PIN disp_val[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END disp_val[4]
  PIN disp_val[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END disp_val[5]
  PIN disp_val[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 847.320 4.000 847.920 ;
    END
  END disp_val[6]
  PIN disp_val[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END disp_val[7]
  PIN disp_val[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1097.560 4.000 1098.160 ;
    END
  END disp_val[8]
  PIN disp_val[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1222.680 4.000 1223.280 ;
    END
  END disp_val[9]
  PIN out_en[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END out_en[0]
  PIN out_en[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.240 4.000 1285.840 ;
    END
  END out_en[10]
  PIN out_en[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1410.360 4.000 1410.960 ;
    END
  END out_en[11]
  PIN out_en[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1535.480 4.000 1536.080 ;
    END
  END out_en[12]
  PIN out_en[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1660.600 4.000 1661.200 ;
    END
  END out_en[13]
  PIN out_en[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2565.970 1756.000 2566.250 1760.000 ;
    END
  END out_en[14]
  PIN out_en[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.090 1756.000 1633.370 1760.000 ;
    END
  END out_en[15]
  PIN out_en[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 1756.000 700.490 1760.000 ;
    END
  END out_en[16]
  PIN out_en[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END out_en[1]
  PIN out_en[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END out_en[2]
  PIN out_en[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END out_en[3]
  PIN out_en[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END out_en[4]
  PIN out_en[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END out_en[5]
  PIN out_en[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END out_en[6]
  PIN out_en[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END out_en[7]
  PIN out_en[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1035.000 4.000 1035.600 ;
    END
  END out_en[8]
  PIN out_en[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1160.120 4.000 1160.720 ;
    END
  END out_en[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2099.530 0.000 2099.810 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 4.670 10.640 2794.040 1749.200 ;
      LAYER met2 ;
        RECT 4.690 1755.720 233.490 1756.000 ;
        RECT 234.330 1755.720 699.930 1756.000 ;
        RECT 700.770 1755.720 1166.370 1756.000 ;
        RECT 1167.210 1755.720 1632.810 1756.000 ;
        RECT 1633.650 1755.720 2099.250 1756.000 ;
        RECT 2100.090 1755.720 2565.690 1756.000 ;
        RECT 2566.530 1755.720 2787.410 1756.000 ;
        RECT 4.690 4.280 2787.410 1755.720 ;
        RECT 4.690 4.000 699.470 4.280 ;
        RECT 700.310 4.000 2099.250 4.280 ;
        RECT 2100.090 4.000 2787.410 4.280 ;
      LAYER met3 ;
        RECT 3.990 1724.160 2787.430 1749.125 ;
        RECT 4.400 1722.760 2787.430 1724.160 ;
        RECT 3.990 1661.600 2787.430 1722.760 ;
        RECT 4.400 1660.200 2787.430 1661.600 ;
        RECT 3.990 1599.040 2787.430 1660.200 ;
        RECT 4.400 1597.640 2787.430 1599.040 ;
        RECT 3.990 1536.480 2787.430 1597.640 ;
        RECT 4.400 1535.080 2787.430 1536.480 ;
        RECT 3.990 1473.920 2787.430 1535.080 ;
        RECT 4.400 1472.520 2787.430 1473.920 ;
        RECT 3.990 1411.360 2787.430 1472.520 ;
        RECT 4.400 1409.960 2787.430 1411.360 ;
        RECT 3.990 1348.800 2787.430 1409.960 ;
        RECT 4.400 1347.400 2787.430 1348.800 ;
        RECT 3.990 1286.240 2787.430 1347.400 ;
        RECT 4.400 1284.840 2787.430 1286.240 ;
        RECT 3.990 1223.680 2787.430 1284.840 ;
        RECT 4.400 1222.280 2787.430 1223.680 ;
        RECT 3.990 1161.120 2787.430 1222.280 ;
        RECT 4.400 1159.720 2787.430 1161.120 ;
        RECT 3.990 1098.560 2787.430 1159.720 ;
        RECT 4.400 1097.160 2787.430 1098.560 ;
        RECT 3.990 1036.000 2787.430 1097.160 ;
        RECT 4.400 1034.600 2787.430 1036.000 ;
        RECT 3.990 973.440 2787.430 1034.600 ;
        RECT 4.400 972.040 2787.430 973.440 ;
        RECT 3.990 910.880 2787.430 972.040 ;
        RECT 4.400 909.480 2787.430 910.880 ;
        RECT 3.990 848.320 2787.430 909.480 ;
        RECT 4.400 846.920 2787.430 848.320 ;
        RECT 3.990 785.760 2787.430 846.920 ;
        RECT 4.400 784.360 2787.430 785.760 ;
        RECT 3.990 723.200 2787.430 784.360 ;
        RECT 4.400 721.800 2787.430 723.200 ;
        RECT 3.990 660.640 2787.430 721.800 ;
        RECT 4.400 659.240 2787.430 660.640 ;
        RECT 3.990 598.080 2787.430 659.240 ;
        RECT 4.400 596.680 2787.430 598.080 ;
        RECT 3.990 535.520 2787.430 596.680 ;
        RECT 4.400 534.120 2787.430 535.520 ;
        RECT 3.990 472.960 2787.430 534.120 ;
        RECT 4.400 471.560 2787.430 472.960 ;
        RECT 3.990 410.400 2787.430 471.560 ;
        RECT 4.400 409.000 2787.430 410.400 ;
        RECT 3.990 347.840 2787.430 409.000 ;
        RECT 4.400 346.440 2787.430 347.840 ;
        RECT 3.990 285.280 2787.430 346.440 ;
        RECT 4.400 283.880 2787.430 285.280 ;
        RECT 3.990 222.720 2787.430 283.880 ;
        RECT 4.400 221.320 2787.430 222.720 ;
        RECT 3.990 160.160 2787.430 221.320 ;
        RECT 4.400 158.760 2787.430 160.160 ;
        RECT 3.990 97.600 2787.430 158.760 ;
        RECT 4.400 96.200 2787.430 97.600 ;
        RECT 3.990 35.040 2787.430 96.200 ;
        RECT 4.400 33.640 2787.430 35.040 ;
        RECT 3.990 10.715 2787.430 33.640 ;
  END
END counter_top
END LIBRARY

